/* Wishbone definitions */

package wb_pkg;
   typedef logic [27:0] adr_t;
   typedef logic [31:0] dat_t;
   typedef logic [3:0]  sel_t;
endpackage

